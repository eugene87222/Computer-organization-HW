//Subject:     CO project 2 - Sign extend
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      楊翔鈞(0516034) 陳柏翰(0516313)
//----------------------------------------------
//Date:        2018/5/2
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module shamt(
    data_i,
    data_o
    );
               
input   [4:0] data_i;
output  [32-1:0] data_o;

reg     [32-1:0] data_o;

always @ ( data_i ) begin
    data_o[31:5] <= 0;
    data_o[4:0] <= data_i[4:0];
  end      
endmodule      
     